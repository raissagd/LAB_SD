sfswfswfsfc